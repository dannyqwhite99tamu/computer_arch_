`timescale 1ns / 1ps
/*
 * Module: InstructionMemory
 *
 * Implements read-only instruction memory
 * 
 */
module InstructionMemory(Data, Address);
   parameter T_rd = 20;
   parameter MemSize = 40;
   
   output [31:0] Data;
   input [63:0]  Address;
   reg [31:0] 	 Data;
   
   /*
    * ECEN 350 Processor Test Functions
    * Texas A&M University
    */
   
   always @ (Address) begin
      #4;
      case(Address)

	/* Test Program 1:
	 * Program loads constants from the data memory. Uses these constants to test
	 * the following instructions: LDUR, ORR, AND, CBZ, ADD, SUB, STUR and B.
	 * 
	 * Assembly code for test:
	 * 
	 * 0: LDUR X9, [XZR, 0x0]    //Load 1 into x9
	 * 4: LDUR X10, [XZR, 0x8]   //Load a into x10
	 * 8: LDUR X11, [XZR, 0x10]  //Load 5 into x11
	 * C: LDUR X12, [XZR, 0x18]  //Load big constant into x12
	 * 10: LDUR X13, [XZR, 0x20]  //load a 0 into X13
	 * 
	 * 14: ORR X10, X10, X11  //Create mask of 0xf
	 * 18: AND X12, X12, X10  //Mask off low order bits of big constant
	 * 
	 * loop:
	 * 1C: CBZ X12, end  //while X12 is not 0
	 * 20: ADD X13, X13, X9  //Increment counter in X13
	 * 24: SUB X12, X12, X9  //Decrement remainder of big constant in X12
	 * 28: B loop  //Repeat till X12 is 0
	 * 2C: STUR X13, [XZR, 0x20]  //store back the counter value into the memory location 0x20
	 */
	

	63'h000: Data = 32'hF84003E9;
	63'h004: Data = 32'hF84083EA;
	63'h008: Data = 32'hF84103EB;
	63'h00c: Data = 32'hF84183EC;
	63'h010: Data = 32'hF84203ED;
	63'h014: Data = 32'hAA0B014A;
	63'h018: Data = 32'h8A0A018C;
	63'h01c: Data = 32'hB400008C;
	63'h020: Data = 32'h8B0901AD;
	63'h024: Data = 32'hCB09018C;
	63'h028: Data = 32'h17FFFFFD;
	63'h02c: Data = 32'hF80203ED;
	63'h030: Data = 32'hF84203ED;  //One last load to place stored value on memdbus for test checking.

	/* *****************Add code for your tests here************* */
	[D29BDE09]->1101||0010||1001||1011||1101||1110||0000||1001|| // MOVZ X9, #0xdef0 LS 0 
	[D2B3578A]->1101||0010||1011||0011||0101||0111||1000||1010|| // MOVZ X10, #0x9abc // LSL16
	[AA09014B]->1010||1010||0000||1001||0000||0001||0100||1011|| // ORR X11, X9, X10 // X11 = 0x000000009abcdef0
	[D2CACF09]->1101||0010||1100||1010||1100||1111||0000||1001|| // MOVZ X9, #0x5678 // LSL32
	[D2E2468A]->1101||0010||1110||0010||0100||0110||1000||1010|| // MOVZ X10, #0x1234 // LSL48
	[AA09014A]->1010||1010||0000||1001||0000||0001||0100||1100|| // ORR X12, X9, X10 // X12 = 0x1234567800000000
	[AA0B0189]->1010||1010||0000||1011||0000||0001||1000||1001|| // ORR  X9, X11, X12 // X9 = 0x123456789abcdef0 
	[8B1F03E0] // ADD X0, XZR, XZR
	[F8028009] // STUR X9, [X0, 0x28]
	[F842800A] // LDUR X10, [X9, 0x28]

			
	default: Data = 32'hXXXXXXXX;
      endcase
   end
endmodule
